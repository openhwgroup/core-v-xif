// Copyright 2024 OpenHW Group.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

module test;

  // eXtension Interface
  /* verilator lint_off UNUSED */
  core_v_xif core_v_xif_bus ();

  initial begin
   $display("Instantiating CORE-V-XIF reference model");
   $finish;
  end

endmodule
